library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity reg12bits is
    port( 
        clk : in std_logic;
        reset : in std_logic;
        wr_en : in std_logic;
        data_in : in signed(11 downto 0);
        data_out : out signed(11 downto 0)
    );
end entity;

architecture a_reg12bits of reg12bits is
    signal registro: signed(11 downto 0) := "000000000000";
begin
    process(clk,reset,wr_en) -- acionado se houver mudança em clk, rst ou wr_en
    begin
        if reset='1' then
            registro <= "000000000000";
        elsif wr_en='1' then
            if rising_edge(clk) then
                registro <= data_in;
            end if;
        end if;
    end process;

    data_out <= registro; -- conexao direta, fora do processo
end architecture;