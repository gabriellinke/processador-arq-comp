library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port( 
        clk : in std_logic;
        address : in unsigned(11 downto 0); -- memória de programa:  1Kbyte = 1024bytes = 4096 bits = 2^12
        data : out unsigned(16 downto 0) := "00000000000000000"
    );
end entity;

architecture a_rom of rom is
    type mem is array (0 to 4095) of unsigned(16 downto 0); -- memória ROM de 1k e com dados de 17 bits (conforme requisitos) - acredito está errado
    constant content_rom : mem := (
        -- caso endereco => conteudo

        -- PROGRAMA LAB 6
        0 => B"01000_011_000000000",  -- LDI R3,000000000B -- P1
        1 => B"01000_100_000000000",  -- LDI R4,000000000B -- P2
        2 => B"00000_100_011_100000", -- ADD R4,R3         -- P3
        3 => B"01000_111_000000001",  -- LDI R7,000000001B -- P4
        4 => B"00000_011_111_100000", -- ADD R4,R3         -- P4
        5 => B"00110_011_000011110",  -- CPI R3,000011110B -- P5
        6 => B"10111_111111111011",   -- BRLO -5           -- P5
        7 => B"00000_101_100_100001", -- MOV R5,R4         -- P6

        -- PROGRAMA PARA TESTAR CP E CPI
        -- 0 => B"01000_001_001100101",  -- LDI R1,001100101B
        -- 1 => B"01000_010_011010011",  -- LDI R2,011010011B
        -- 2 => B"00000_001_010_100110", -- CP  R1,R2
        -- 3 => B"00110_001_000000001",  -- CPI R1,000000001B
        -- 4 => B"00110_001_011111111",  -- CPI R1,011111111B
        -- 5 => B"00110_001_001100101",  -- CPI R1,001100101B
        -- 6 => B"00110_010_000000001",  -- CPI R2,000000001B
        -- 7 => B"00110_010_011111111",  -- CPI R2,011111111B
        -- 8 => B"00110_010_011010011",  -- CPI R2,011010011B
        -- 9 => B"00000_001_000_100000", -- ADD R1,R0
        -- 10 => B"00000_010_000_100000", -- ADD R2,R0

        -- PROGRAMA LAB 5
        -- 0 => B"01000_011_000000101",    -- LDI R3,000000101B
        -- 1 => B"01000_100_000001000",    -- LDI R4,000001000B
        -- 2 => B"00000_011_100_100000",   -- ADD R3,R4
        -- 3 => B"00000_101_011_100001",   -- MOV R5,R3
        -- 4 => B"00010_101_000000001",    -- SUBI R1,000000001B
        -- 5 => B"11111_000000010100",     -- JMP 20
        -- 20 => B"00000_011_101_100001",  -- MOV R3,R5
        -- 21 => B"11111_000000000010",    -- JMP 2

        -- PROGRAMA PARA TESTAR AS INSTRUCOES BASICAS
        -- 0 => B"01000_001_000000100", -- LDI 001 000000100
        -- 1 => B"01000_001_010000000", -- LDI 001 010000000
        -- 2 => B"01000_010_000000001", -- LDI 010 000000001
        -- 3 => B"00010_001_000000001", --SUBI 001 000000001
        -- 4 => B"00010_010_000000100", --SUBI 010 000000100
        -- 5 => B"00000_001_000_100000", -- ADD 001 000
        -- 6 => B"01000_111_000001100", -- LDI 111 000001100
        -- 7 => B"01000_110_010010001", -- LDI 110 010010001
        -- 8 => B"00000_111_110_100000", -- ADD 111 110
        -- 9 => B"00000_111_110_100010", -- SUB 111 110
        -- 10 => B"00000_111_001_100001", -- MOV 111 001
        -- 11 => B"00000_110_010_100001", -- MOV 110 001
        -- 12 => B"00000_111_000_100000", -- ADD 111 000
        -- 13 => B"00000_110_000_100000", -- ADD 110 000
        -- 14 => B"11111_000000000000", -- jump para 0

        -- 0 => "11111000000000111", -- jump para 7
        -- 1 => "00001010110110000",
        -- 2 => "00000000000011111",
        -- 3 => "11111000000000101", -- jump para 5
        -- 4 => "11111000000001000", -- jump para 8
        -- 5 => "00000000001111110",
        -- 6 => "11111000000000100", -- jump para 4
        -- 7 => "11111000000000001", -- jump para 1
        -- 8 => "00000001100001001",
        -- 9 => "11100000000001010",
        -- 10 => "00011000000001011",
        -- 11 => B"00010_001_000000001", --SUBI 001 000000001
        -- 12 => B"00010_001_000000100", --SUBI 001 000000100
        -- 13 => B"00010_010_000000010", --SUBI 010 000000010
        -- 14 => B"00000_001_010_100000", -- ADD 001 010
        -- abaixo: casos omissos => (zero em todos os bits)
        others => (others=>'0')
    );
begin
    process(clk)
    begin
        if(rising_edge(clk)) then
            data <= content_rom(to_integer(address));
        end if;
    end process;
end architecture;