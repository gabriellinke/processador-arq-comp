library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port( 
        clk : in std_logic;
        address : in unsigned(11 downto 0); -- memória de programa:  1Kbyte = 1024bytes = 4096 bits = 2^12
        data : out unsigned(16 downto 0) := "00000000000000000"
    );
end entity;

architecture a_rom of rom is
    type mem is array (0 to 4095) of unsigned(16 downto 0); -- memória ROM de 1k e com dados de 17 bits (conforme requisitos) - acredito está errado
    constant content_rom : mem := (
        -- caso endereco => conteudo    

        -- PROGRAMA DE VALIDACAO
        -- loop para preencher quantidade especificada de numeros
        0 => B"01000_110_000100000",    -- LDI R6,32 -- número limite
		1 => B"01000_001_000000000",    -- LDI R1,0
		2 => B"01000_111_000000000",    -- LDI R7,0
		3 => B"00010_001_111111111",    -- SUBI R1,-1
		4 => B"00010_111_111111111",    -- SUBI R7,-1
		5 => B"01101_001_000000000",    -- ST R1
		6 => B"00000_001_110_100110",   -- CP R7,R6
		7 => B"10111_111111111011",     -- BRLO -5  

        -- loop para remover os nao primos
        8 => B"01000_010_000000001",    -- LDI R2,1
		9 => B"01000_111_000000000",    -- LDI R7,0
		10 => B"00010_010_111111111",   -- SUBI R2,-1
		11 => B"00000_111_010_100000",  -- ADD R7,R2
		12 => B"01100_100_000000000",   -- LD R4
        13 => B"00000_100_000_100110",  -- CP R4,R0
        14 => B"10100_000000000100",    -- BREQ 4
		15 => B"00000_111_100_100000",  -- ADD R7,R4
		16 => B"01101_000_000000000",   -- ST R0
		17 => B"00000_111_110_100110",  -- CP R7,R6
		18 => B"10111_111111111100",    -- BRLO -4

		19 => B"00000_010_110_100110",  -- CP R2,R6
		20 => B"10111_111111110100",    -- BRLO -12

        -- loop para ler a memoria do 2 ao 32
        21 => B"01000_111_000000001",   -- LDI R7,1
		22 => B"00010_111_111111111",   -- SUBI R7,-1
		23 => B"01100_011_000000000",   -- LD R3
		24 => B"00000_111_110_100110",  -- CP R7,R6
		25 => B"10111_111111111100",    -- BRLO -4
        -- FIM DO PROGRAMA DE VALIDACAO 

        -- PROGRAMA PARA TESTAR LD E ST
        -- Testa se os dados estão ficando salvos na memória e se os valores nos registradores não estão sendo sobrescritos em nenhum momento
        -- 0 => B"01000_001_000000101",   --  LDI R1,000000101B -- 5
        -- 1 => B"01000_010_011111111",   --  LDI R2,011111111B -- 255
        -- 2 => B"01000_011_000000000",   --  LDI R3,000000000B -- 0
        -- 3 => B"01000_100_010110100",   --  LDI R4,010110100B -- 180
        -- 4 => B"01000_101_010001111",   --  LDI R5,010001111B -- 143
        -- 5 => B"01000_110_000000001",   --  LDI R6,000000001B -- 1

        -- 6 => B"01000_111_000000000",   --  LDI R7,000000000B -- 0
        -- 7 => B"01101_001_000000000",   --  ST R1
        -- 8 => B"01000_111_001010111",   --  LDI R7,001010111B -- 87
        -- 9 => B"01101_010_000000000",   --  ST R2
        -- 10 => B"01000_111_000101010",  --  LDI R7,000101010B -- 42
        -- 11 => B"01101_011_000000000",  --  ST R3
        -- 12 => B"01000_111_000010011",  --  LDI R7,000010011B -- 19
        -- 13 => B"01101_100_000000000",  --  ST R4
        -- 14 => B"01000_111_001111111",  --  LDI R7,001111111B -- 127
        -- 15 => B"01101_101_000000000",  --  ST R5
        -- 16 => B"01000_111_001100100",  --  LDI R7,001100100B -- 100
        -- 17 => B"01101_110_000000000",  --  ST R6

        -- 18 => B"00000_001_000_100000", --  ADD R1,R0
        -- 19 => B"01000_111_000000000",  --  LDI R7,000000000B -- 0
        -- 20 => B"01100_001_000000000",  --  LD R1
        -- 21 => B"00000_001_000_100000", --  ADD R1,R0
         
        -- 22 => B"01000_111_001010111",  --  LDI R7,001010111B -- 87
        -- 23 => B"01100_001_000000000",  --  LD R1
        -- 24 => B"00000_001_010_100000", --  ADD R1,R2

        -- 25 => B"01000_111_000101010",  --  LDI R7,000101010B -- 42
        -- 26 => B"01100_001_000000000",  --  LD R1
        -- 27 => B"00000_001_011_100000", --  ADD R1,R3

        -- 28 => B"01000_111_000010011",  --  LDI R7,000010011B -- 19
        -- 29 => B"01100_001_000000000",  --  LD R1
        -- 30 => B"00000_001_100_100000", --  ADD R1,R4

        -- 31 => B"01000_111_001111111",  --  LDI R7,001111111B -- 127
        -- 32 => B"01100_001_000000000",  --  LD R1
        -- 33 => B"00000_001_101_100000", --  ADD R1,R5

        -- 34 => B"01000_111_001100100",  --  LDI R7,001100100B -- 100
        -- 35 => B"01100_001_000000000",  --  LD R1
        -- 36 => B"00000_001_110_100000", --  ADD R1,R6

        -- --Testa se a memória consegue armazenar valores maiores (Deixar o 16º bit como 1)
        -- 37 => B"01000_110_111111110",  --  LDI R6,111111110B -- -2
        -- 38 => B"01000_111_000010000",  --  LDI R7,000010000B -- 16
        -- 39 => B"01101_110_000000000",  --  ST R6
        -- 40 => B"01100_010_000000000",  --  LD R2
        -- 41 => B"01000_110_000010010",  --  LDI R6,000010010B -- 18
        -- 42 => B"00000_110_010_100000", --  ADD R6,R2
        
        -- -- Lê um endereço que não foi utilizado para ver se retorna undefined
        -- 43 => B"01000_111_000000001",  --  LDI R7,000000001B -- 1
        -- 44 => B"01100_010_000000000",  --  LD R2

        -- -- Testa se é possível reescrever num mesmo endereço de memória. Também testa nova escrita no endereço ao lado.
        -- 45 => B"01000_111_000000000",  --  LDI R7,000000000B -- 0
        -- 46 => B"01000_001_111110001",  --  LDI R1,111110001B -- -15
        -- 47 => B"01101_001_000000000",  --  ST R1
        -- 48 => B"01000_001_000001101",  --  LDI R1,000001101B -- 13
        -- 49 => B"00010_111_111111111",  --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 50 => B"01101_001_000000000",  --  ST R1

        -- 51 => B"01000_111_001010111",  --  LDI R7,001010111B -- 87
        -- 52 => B"01000_010_101011011",  --  LDI R2,101011011B -- -165
        -- 53 => B"01101_010_000000000",  --  ST R2
        -- 54 => B"01000_010_000011010",  --  LDI R2,000001101B -- 26
        -- 55 => B"00010_111_111111111",  --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 56 => B"01101_010_000000000",  --  ST R2

        -- 57 => B"01000_111_000101010",  --  LDI R7,000101010B -- 42
        -- 58 => B"01000_011_111011011",  --  LDI R3,111011011B -- -37
        -- 59 => B"01101_011_000000000",  --  ST R3
        -- 60 => B"01000_011_000000110",  --  LDI R3,000000110B -- 6
        -- 61 => B"00010_111_111111111",  --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 62 => B"01101_011_000000000",  --  ST R3

        -- 63 => B"01000_111_000010011",  --  LDI R7,000010011B -- 19
        -- 64 => B"01000_100_111111110",  --  LDI R4,111111110B -- -2
        -- 65 => B"01101_100_000000000",  --  ST R4
        -- 66 => B"01000_100_000000000",  --  LDI R4,000000000B -- 0
        -- 67 => B"00010_111_111111111",  --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 68 => B"01101_100_000000000",  --  ST R4

        -- 69 => B"01000_111_001111111",  --  LDI R7,001111111B -- 127
        -- 70 => B"01000_101_110101001",  --  LDI R5,110101001B -- -87
        -- 71 => B"01101_101_000000000",  --  ST R5
        -- 72 => B"01000_101_000001001",  --  LDI R5,000001001B -- 9
        -- 73 => B"00010_111_111111111",  --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 74 => B"00000000000000000",    --  NOP                     - Como a memória só vai até 127, se tentar gravar no 128 vai acabar gravando por cima do que tem no 0

        -- 75 => B"01000_111_001100100",  --  LDI R7,001100100B -- 100
        -- 76 => B"01000_110_111011000",  --  LDI R6,111011000B -- -40
        -- 77 => B"01101_110_000000000",  --  ST R6
        -- 78 => B"01000_110_000000100",  --  LDI R6,000000100B -- 4
        -- 79 => B"00010_111_111111111",  --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 80 => B"01101_110_000000000",  --  ST R6
        
        -- -- Carrega os valores salvos em memória em diferentes registradores, pra ver se é possível usar o LD em todos eles.
        -- 81 => B"01000_111_000000000",  --  LDI R7,000000000B -- 0
        -- 82 => B"01100_011_000000000",  --  LD R3
        -- 83 => B"00010_111_111111111",  --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 84 => B"01100_101_000000000",  --  LD R5
        -- 85 => B"00000_011_101_100000", --  ADD R3,R5

        -- 86 => B"01000_111_001010111",  --  LDI R7,001010111B -- 87
        -- 87 => B"01100_001_000000000",  --  LD R1
        -- 88 => B"00010_111_111111111",  --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 89 => B"01100_010_000000000",  --  LD R4
        -- 90 => B"00000_001_010_100000", --  ADD R1,R4

        -- 91 => B"01000_111_000101010",  --  LDI R7,000101010B -- 42
        -- 92 => B"01100_010_000000000",  --  LD R2
        -- 93 => B"00010_111_111111111",  --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 94 => B"01100_110_000000000",  --  LD R6
        -- 95 => B"00000_010_110_100000", --  ADD R2,R6

        -- 96 => B"01000_111_000010011",  --  LDI R7,000010011B -- 19
        -- 97 => B"01100_010_000000000",  --  LD R2
        -- 98 => B"00010_111_111111111",  --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 99 => B"01100_001_000000000",  --  LD R1
        -- 100 => B"00000_001_010_100000",--  ADD R1,R2

        -- 101 => B"01000_111_001111111", --  LDI R7,001111111B -- 127
        -- 102 => B"01100_110_000000000", --  LD R6
        -- 103 => B"00000_001_110_100000",--  ADD R1,R6

        -- 104 => B"01000_111_001100100", --  LDI R7,001100100B -- 100
        -- 105 => B"01100_010_000000000", --  LD R4
        -- 106 => B"00010_111_111111111", --  SUBI R7,111111111B-- -1 - faz o mesmo que faria um ADDI R7,1
        -- 107 => B"01100_101_000000000", --  LD R5
        -- 108 => B"00000_010_101_100000",--  ADD R4,R5

        -- Programa de teste com branches
        -- let a = 0;

        -- for(let i=0; i<30; i++)
        --     a+=1;
        
        -- if(a==30)
        --     a+=5;
        -- else
        --     a-=5
        --
        -- for(let i=25; i>=1; i--)
        --     a-=1;
        
        -- if(a!=0)
        --     a+=100
        -- else
        --     a-=100        

        -- 0 => B"01000_001_000000000",  --LDI R1,000000000B
        -- 1 => B"01000_110_000000000",  --LDI R6,000000000B
        -- 2 => B"01000_111_000000001",  --LDI R7,000000001B
        -- 3 => B"00000_001_111_100000", --ADD R1,R7
        -- 4 => B"00000_110_111_100000", --ADD R6,R7
        -- 5 => B"00110_110_000011110",  --CPI R6,000011110B
        -- 6 => B"10111_111111111100",   --BRLO -4
        -- 7 => B"00110_001_000011110",  --CPI R1,000011110B
        -- 8 => B"10101_000000000011",   --BRNE 3
        -- 9 => B"01000_101_000000101",  --LDI R5,000000101B
        -- 10 => B"00000_001_101_100000",--ADD R1,R5
        -- 11 => B"10000_000000000001",  --RJMP 1
        -- 12 => B"00010_001_000000101", --SUBI R1,000000101B

        -- 13 => B"01000_110_000011001", --LDI R6,000011001B
        -- 14 => B"00010_001_000000001", --SUBI R1,000000001B
        -- 15 => B"00010_110_000000001", --SUBI R6,000000001B
        -- 16 => B"00110_110_000000001", --CPI R6,000000001B
        -- 17 => B"10110_111111111100",  --BRSH -4

        -- 18 => B"00110_001_000000000", --CPI R1,000000000B
        -- 19 => B"10100_000000000011",  --BREQ 3
        -- 20 => B"01000_101_001100100", --LDI R5,001100100B
        -- 21 => B"00000_001_101_100000",--ADD R1,R5
        -- 22 => B"10000_000000000001",  --RJMP 1
        -- 23 => B"00010_001_001100100", --SUBI R1,001100100B

        -- PROGRAMA LAB 6
        -- 0 => B"01000_011_000000000",  -- LDI R3,000000000B -- P1
        -- 1 => B"01000_100_000000000",  -- LDI R4,000000000B -- P2
        -- 2 => B"00000_100_011_100000", -- ADD R4,R3         -- P3
        -- 3 => B"01000_111_000000001",  -- LDI R7,000000001B -- P4
        -- 4 => B"00000_011_111_100000", -- ADD R4,R3         -- P4
        -- 5 => B"00110_011_000011110",  -- CPI R3,000011110B -- P5
        -- 6 => B"10111_111111111011",   -- BRLO -5           -- P5
        -- 7 => B"00000_101_100_100001", -- MOV R5,R4         -- P6

        -- PROGRAMA PARA TESTAR CP E CPI
        -- 0 => B"01000_001_001100101",  -- LDI R1,001100101B
        -- 1 => B"01000_010_011010011",  -- LDI R2,011010011B
        -- 2 => B"00000_001_010_100110", -- CP  R1,R2
        -- 3 => B"00110_001_000000001",  -- CPI R1,000000001B
        -- 4 => B"00110_001_011111111",  -- CPI R1,011111111B
        -- 5 => B"00110_001_001100101",  -- CPI R1,001100101B
        -- 6 => B"00110_010_000000001",  -- CPI R2,000000001B
        -- 7 => B"00110_010_011111111",  -- CPI R2,011111111B
        -- 8 => B"00110_010_011010011",  -- CPI R2,011010011B
        -- 9 => B"00000_001_000_100000", -- ADD R1,R0
        -- 10 => B"00000_010_000_100000", -- ADD R2,R0

        -- PROGRAMA LAB 5
        -- 0 => B"01000_011_000000101",    -- LDI R3,000000101B
        -- 1 => B"01000_100_000001000",    -- LDI R4,000001000B
        -- 2 => B"00000_011_100_100000",   -- ADD R3,R4
        -- 3 => B"00000_101_011_100001",   -- MOV R5,R3
        -- 4 => B"00010_101_000000001",    -- SUBI R1,000000001B
        -- 5 => B"11111_000000010100",     -- JMP 20
        -- 20 => B"00000_011_101_100001",  -- MOV R3,R5
        -- 21 => B"11111_000000000010",    -- JMP 2

        -- PROGRAMA PARA TESTAR AS INSTRUCOES BASICAS
        -- 0 => B"01000_001_000000100", -- LDI 001 000000100
        -- 1 => B"01000_001_010000000", -- LDI 001 010000000
        -- 2 => B"01000_010_000000001", -- LDI 010 000000001
        -- 3 => B"00010_001_000000001", --SUBI 001 000000001
        -- 4 => B"00010_010_000000100", --SUBI 010 000000100
        -- 5 => B"00000_001_000_100000", -- ADD 001 000
        -- 6 => B"01000_111_000001100", -- LDI 111 000001100
        -- 7 => B"01000_110_010010001", -- LDI 110 010010001
        -- 8 => B"00000_111_110_100000", -- ADD 111 110
        -- 9 => B"00000_111_110_100010", -- SUB 111 110
        -- 10 => B"00000_111_001_100001", -- MOV 111 001
        -- 11 => B"00000_110_010_100001", -- MOV 110 001
        -- 12 => B"00000_111_000_100000", -- ADD 111 000
        -- 13 => B"00000_110_000_100000", -- ADD 110 000
        -- 14 => B"11111_000000000000", -- jump para 0

        -- PROGRAMA PARA TESTAR AS INSTRUCOES DE BRANCH
        -- 1 => B"01000_010_000000001", -- LDI R2,000000001B
        -- 2 => B"01000_001_000000000", -- LDI R1,000000000B
        -- 3 => B"00000_001_010_100000", -- ADD R1,R2
        -- 4 => B"00110_001_000000010", -- CPI R1,000000010B
        -- 11 => B"10100_111111111101", -- BREQ -3
        -- 12 => B"01000_001_000000000", -- LDI R1,000000000B
        -- 13 => B"00000_001_010_100000", -- ADD R1,R2
        -- 14 => B"00110_001_000000001", -- CPI R1,000000001B
        -- 15 => B"10101_111111111101", -- BRNE -3
        -- 16 => B"01000_001_000000111", -- LDI R1,000000111B
        -- 17 => B"00000_001_010_100010", -- SUB R1,R2
        -- 18 => B"00110_001_000000001", -- CPI R1,000000001B
        -- 19 => B"10110_111111111101", -- BRSH -3
        -- 20 => B"01000_001_000000000", -- LDI R1,000000000B
        -- 21 => B"00000_001_010_100000", -- ADD R1,R2
        -- 22 => B"00110_001_000000110", -- CPI R1,000000001B
        -- 23 => B"10111_111111111101", -- BRLO -3

        -- 0 => "11111000000000111", -- jump para 7
        -- 1 => "00001010110110000",
        -- 2 => "00000000000011111",
        -- 3 => "11111000000000101", -- jump para 5
        -- 4 => "11111000000001000", -- jump para 8
        -- 5 => "00000000001111110",
        -- 6 => "11111000000000100", -- jump para 4
        -- 7 => "11111000000000001", -- jump para 1
        -- 8 => "00000001100001001",
        -- 9 => "11100000000001010",
        -- 10 => "00011000000001011",
        -- 11 => B"00010_001_000000001", --SUBI 001 000000001
        -- 12 => B"00010_001_000000100", --SUBI 001 000000100
        -- 13 => B"00010_010_000000010", --SUBI 010 000000010
        -- 14 => B"00000_001_010_100000", -- ADD 001 010
        -- abaixo: casos omissos => (zero em todos os bits)
        others => (others=>'0')
    );
begin
    process(clk)
    begin
        if(rising_edge(clk)) then
            data <= content_rom(to_integer(address));
        end if;
    end process;
end architecture;